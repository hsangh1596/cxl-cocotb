module CMSS_TOP_WRAPPER
   ()
   ;
endmodule
